module surrogate_engine():
endmodule
