

`timescale 1ns/1ps

module tb_top_snn1();

//////////////////////////////////////////////////////////////
// Signals
//////////////////////////////////////////////////////////////

reg clk;
reg rst;
reg start;
wire done;

//////////////////////////////////////////////////////////////
// DUT
//////////////////////////////////////////////////////////////

top_snn uut (
    .clk(clk),
    .rst(rst),
    .start(start),
    .done(done)
);

//////////////////////////////////////////////////////////////
// Clock Generation (100 MHz)
//////////////////////////////////////////////////////////////

initial begin
    clk = 0;
    forever #5 clk = ~clk;   // 10ns period
end

//////////////////////////////////////////////////////////////
// Reset + Start Sequence
//////////////////////////////////////////////////////////////

initial begin
    rst = 1;
    start = 0;

    // Hold reset for 20ns
    #20;
    rst = 0;

    // Wait 20ns
    #20;

    // Give start pulse
    start = 1;
    #10;
    start = 0;

    // Wait long enough for full computation
    #5000;

    $finish;
end

//////////////////////////////////////////////////////////////
// Monitor
//////////////////////////////////////////////////////////////

initial begin
    $monitor("Time=%0t | state=%0d | neuron=%0d | input=%0d | acc=%0d | done=%b",
              $time,
              uut.state,
              uut.neuron_idx,
              uut.input_idx,
              uut.accumulator,
              done);
end

endmodule
