`timescale 1ns/1ps

module tb_mem_controller;

reg clk;
reg we;
reg [15:0] addr;
reg [31:0] wdata;
wire [31:0] rdata;

//////////////////////////////////////////////////////////////
// DUT
//////////////////////////////////////////////////////////////

snn_mem_controller uut (
    .clk(clk),
    .we(we),
    .addr(addr),
    .wdata(wdata),
    .rdata(rdata)
);

//////////////////////////////////////////////////////////////
// Clock
//////////////////////////////////////////////////////////////

always #5 clk = ~clk;

//////////////////////////////////////////////////////////////
// Test Sequence
//////////////////////////////////////////////////////////////

initial begin
    clk = 0;
    we  = 0;
    addr = 0;
    wdata = 0;

    //////////////////////////////////////////////////////////
    // TEST BANK0 (0x0000)
    //////////////////////////////////////////////////////////
    #10;
    addr  = 16'h0000;
    wdata = 32'hDEADBEEF;
    we    = 1;
    #10;
    we    = 0;

    #10;
    addr  = 16'h0000;
    #10;

    //////////////////////////////////////////////////////////
    // TEST BANK1 (0x1000)
    //////////////////////////////////////////////////////////
    addr  = 16'h1000;
    wdata = 32'h11112222;
    we    = 1;
    #10;
    we    = 0;

    #10;
    addr = 16'h1000;
    #10;

    //////////////////////////////////////////////////////////
    // TEST BANK3 (0x4000)
    //////////////////////////////////////////////////////////
    addr  = 16'h4000;
    wdata = 32'h33334444;
    we    = 1;
    #10;
    we    = 0;

    #10;
    addr = 16'h4000;
    #10;

    //////////////////////////////////////////////////////////
    // TEST BANK5 (0xE000)
    //////////////////////////////////////////////////////////
    addr  = 16'hE000;
    wdata = 32'hAAAA5555;
    we    = 1;
    #10;
    we    = 0;

    #10;
    addr = 16'hE000;
    #10;

    $stop;
end

endmodule
