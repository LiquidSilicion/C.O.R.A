`timescale 1ns / 1ps

module tb_top_snn;

//////////////////////////////////////////////////////////////
// Testbench Signals
//////////////////////////////////////////////////////////////

reg clk;
reg rst;
reg start;
wire done;

//////////////////////////////////////////////////////////////
// Instantiate DUT
//////////////////////////////////////////////////////////////

top_snn uut (
    .clk(clk),
    .rst(rst),
    .start(start),
    .done(done)
);

//////////////////////////////////////////////////////////////
// Clock Generation (10ns period = 100MHz)
//////////////////////////////////////////////////////////////

initial begin
    clk = 0;
    forever #5 clk = ~clk;
end

//////////////////////////////////////////////////////////////
// Stimulus
//////////////////////////////////////////////////////////////

initial begin

    // Initialize
    rst   = 1;
    start = 0;

    // Hold reset
    #50;
    rst = 0;

    // Wait a little
    #20;

    // Pulse start for 1 cycle
    start = 1;
    #10;
    start = 0;

    // Wait for done
    wait(done);

    #50;

    $stop;
end

endmodule
