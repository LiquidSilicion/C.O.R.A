module input_from_aer();
  input clk,
  input rst_n,
  input wire [31:0]in,
  input aer_valid,
  
  
  output reg [3:0]channel_Id,
  output reg [23:0]timestamp;
  
  always@


endmodule
